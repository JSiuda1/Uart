module uart_rx(
	input clk,
	input rx,
);